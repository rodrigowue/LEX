.subckt AN4D8BWP16P90CPD A1 A2 A3 A4 Z VDD VSS VPP VBB
XMM16_1 net26 A3 VDD VPP P12 L=0.016u nfin=4 as=5.698e-15
XMM16_2 net26 A3 VDD VPP P12 L=0.016u nfin=4
XMM16_3 net26 A3 VDD VPP P12 L=0.016u nfin=4 as=5.698e-15
XMM17_1 net26 A1 VDD VPP P12 L=0.016u nfin=4 as=5.544e-15
XMM17_2 net26 A1 VDD VPP P12 L=0.016u nfin=4
XMM17_3 net26 A1 VDD VPP P12 L=0.016u nfin=4 as=5.698e-15
XMM18_1 net26 A2 VDD VPP P12 L=0.016u nfin=4
XMM18_2 net26 A2 VDD VPP P12 L=0.016u nfin=4 as=5.698e-15
XMM18_3 net26 A2 VDD VPP P12 L=0.016u nfin=4
XMM19_1 net030 A2 net034 VBB N12 L=0.016u nfin=4
XMM19_2 net030 A2 net034 VBB N12 L=0.016u nfin=4 as=5.698e-15
XMM19_3 net030 A2 net034 VBB N12 L=0.016u nfin=4
XMM20_1 net034 A3 net038 VBB N12 L=0.016u nfin=4
XMM20_2 net034 A3 net038 VBB N12 L=0.016u nfin=4 as=5.698e-15
XMM20_3 net034 A3 net038 VBB N12
XMM21_1 net038 A4 VSS VBB N12 L=0.016u nfin=4
XMM21_2 net038 A4 VSS VBB N12 L=0.016u nfin=4 as=5.698e-15
XMM21_3 net038 A4 VSS VBB N12 L=0.016u nfin=4
XMM22_1 net26 A1 net030 VBB N12 L=0.016u nfin=4
XMM22_2 net26 A1 net030 VBB N12 L=0.016u nfin=4 as=5.698e-15
XMM22_3 net26 A1 net030 VBB N12 L=0.016u nfin=4
XMM23_1 net26 A4 VDD VPP P12 L=0.016u nfin=4
XMM23_2 net26 A4 VDD VPP P12 L=0.016u nfin
XMM23_3 net26 A4 VDD VPP P12 L=0.016u nfin=4
XMM4_1 Z net26 VDD VPP P12 L=0.016u nfin=4 as=5.698e-15
XMM4_2 Z net26 VDD VPP P12 L=0.016u nfin=4
XMM4_3 Z net26 VDD VPP P12 L=0.016u nfin=4 as=5.698e-15
XMM4_4 Z net26 VDD VPP P12 L=0.016u nfin=4
XMM4_5 Z net26 VDD VPP P12 L=0.016u nfin=4 as=5.698e-15
XMM4_6 Z net26 VDD VPP P12 L=0.016u nfin=4
XMM4_7 Z net26 VDD VPP P12
XMM4_8 Z net26 VDD VPP P12 L=0.016u nfin=4
XMM5_1 Z net26 VSS VBB N12 L=0.016u nfin=4 as=5.698e-15
XMM5_2 Z net26 VSS VBB N12 L=0.016u nfin=4
XMM5_3 Z net26 VSS VBB N12 L=0.016u nfin=4 as=5.698e-15
XMM5_4 Z net26 VSS VBB N12 L=0.016u nfin=4
XMM5_5 Z net26 VSS VBB N12 L=0.016u nfin=4 as=5.698e-15
XMM5_6 Z net26 VSS VBB N12 L=0.016u nfin=4
XMM5_7 Z net26 VSS VBB N12 L=0.016u nfin=4 as=5.698e-15
XMM5_8 Z net26 VSS VBB N12 L=0.016u nfin=4
.ends
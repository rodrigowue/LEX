.subckt sky130_fd_sc_hs__buf_1 A VGND VNB VPB VPWR X
X0 VGND a_27_164# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_27_164# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X2 a_27_164# A VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X3 VPWR a_27_164# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
.ends
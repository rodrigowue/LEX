.SUBCKT NAND3D0BWP A B C OUT VDD VSS
*.pininfo A:I B:I C:I OUT:O VSS:G VDD:P
MP0 VDD A OUT VDD PCH W=2.5E-06 L=0.04E-06
MP1 VDD B OUT VDD PCH W=2.5E-06 L=0.04E-06
MP2 VDD C OUT VDD PCH W=2.5E-06 L=0.04E-06
MN0 OUT A rand0 VSS NCH W=2.5E-06 L=0.04E-06
MN1 rand0 B rand1 VSS NCH W=2.5E-06 L=0.04E-06
MN2 rand1 C VSS VSS NCH W=2.5E-06 L=0.04E-06

.ENDS


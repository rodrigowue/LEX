.subckt sky130_fd_sc_hs__xnor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_376_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X1 a_293_74# a_138_385# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_112_119# B a_138_385# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VGND B a_293_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VGND A a_112_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 VPWR A a_138_385# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X6 a_293_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_138_385# B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X8 a_376_368# B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
X9 Y a_138_385# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=150000u
.ends